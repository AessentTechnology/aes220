x�\��,���(�������G%n���-;�ml%($E% ���kϴ��ɶu�+�w�+�����7�m��\!;	�����kE��KE����m߸�mDmc�F �$Ab�4��C�?�)67�+���7�-��M��L	�����]Ce�]K�ջ�-ի�mE,�D%!����5��6?�+�)����Ȇ]`D\�� `�����GI��CEl��m�{0aD�*�De�lOkƵ����u*�w�)�?���8�l%x�\	��$���M-/�Cn׻�mo��mE%(�d)����4�ꉤe�/�5�+5�������\��Xˉ�	���CD�=CM����o׺�mDW`�DE 4ajäA��&g�o�V�*5���5p|��Ta����B�Ce��c�G��m�s�-D`�!�������ôw#6u�+׽������V!��v����ߩ-�MGE��CE斻4,W��dD �L0����ʴ�胶w5+�wu"���5%����_z|�TA���B�i���ce��cef��	eǱ�mD �d%!�������c�vuk�w�)��1u��6�\!xn|��������e��cElU� -ǫ�md(D$����O���˶w-�7+���=7�&\!x�L	� ��	%��Ce�}!���-ջm@a�DE@�,ꧬ�*�?w�+�'�+���5����|	��L	���ʛ���}%E��ae.W��m���m ���I��AjA5�+��+���5��h�L��\���B�	���	E��GE�W=�-׻�mE!�d(4�j˴A�C�g�)?�/�������|	�\������ ��Ce��M%�-���m!� �5��s��j�&w�+�7#����řU��~!چt���ï�"��Ca��CE�׿�mӲ�}d�d �p���$���vr;�v�#��g�����\��u!�	j�;��B�SE��SEf���lS��mD
(�Cj�4@��u�+�u�#���3ݽ9�'ie�#�~M��,l��MK,�uQg�tgG��EFM2QBt&,Q���l!��ud0�b�fAa�'HG�'��l�$N6�v�Av�o���gG��G;}BE2UjG.$�G<���t!��T!��Yb��g�e�#Y$�/=4l��4l�!v�.�2�gg��'W=xEpUBE25FQ/lEn'���r#��u ��d��bIa�'Ie�!�<l��<h�f"�.�v`k��gO�|@3BEcUb}.lE&�mtA��t%d��Gt�FIe�Iw�7�<l��<h�n�nI�w�e�]|g���U2UBEbuBo�U.m�tA��`a��D���vIE�DMe�'/4O4�h�
v�v�cc��F�uE>qBE6UBU.�U.E��|!��tapϙfuW��ae�#Ie�&�<`t�<l�.�vH�v�g�?�g��2 M"eBu/�U.���t!��d!�m�o�dIe{'I}�'�<d$�<e��f�v�bG�gƏ�dUBm3EB.mQ.��eta��t!��jp�fK%-I`�'�<d0�<lt\�t�V�t�cǟ�w�/�G2uG%s]bUWA�u.���t#�at!�	fQ�n�e�%aE�%<l�� I�
�fLV�gş�f��f6UBG2TFu.�E.$�mt0�61���f�fI-}e�-�-l�,l�.	��dIg���e���M2Ug2U].�U/%��4!��t!���o��lIm�'Ie?'�=-��=l4w��v�e�tgg��e"uBe0]BE/�U$���p!�yt!��dt��gIe�gIeo'�ul��|h�Pf��v�kG�w��e"]BErEbT>�Un%n��|a��p#�gt��mAe�*Aa�&(l �~m��&h.rIwd��g��g2uR2CQ.!�.̏�t1W�$!���&~��teogke�'�<h��<|��r��V�gǟyg׏�E X@A&uBu.lU,h��t!��ta��v��f�E�gHe�'�<l��4$4�u�,�b���i!��!!w_f�-tn6��Ѽ��qg5�&/RhoO�H|��N�����'+0�&82�oKM	nEo0|\��_VbQBLQ؉!Q�� gg�	�$�+�M~�M~��n�����&+�#_KO_I)kO�Ry�VL�XRLY@G�ҡ!���!nE��g�)Dx�D>��S��nqg{+�'?2�%O	oNM�tT��VX�	bOQbMUЍ)�Qi#�'r
�e��M~	]>�7쓼?.�%|�%o�oO-)kJ	>\��F\�[PLy;Bd��i��!gw�gvAMn�KM{����+���'��7oho_	n	�FT֞_\�hbLr�а QP�!�gu*�gWO�JM	KM~���Ӿ��SwDJ"=2�+O	kf-I>V\m�VT�x?cFYj\Q�	!aP�!kf�#u��i~�Km~����=��'?2j#/#�`G!oOI	�Vt��V]�]_B\IBL��)!��[a�g�+�KWK�M^�	O~"��Ӿ���'Y�'?J/oy+c	�V\��VT�JBLYRL�P�!�Ҁc�d��g�C�M~�E~*�3>���'~Cjs?��O@oNMm�Rt��fS�]~`LX?b|�ө �p�!57�	vuK�L~�kol��fӮ�f�'?A'6�gOi_	�\|�v�Y/@,y_jLQЈ!��H!�g�	�%v)i~�od>�jS>���'?�&?ފnOl[M	]D\��F\-QRLX6L���)��-�gugw+
M:!)~�3�Ӯ�n�g?R�'?IOOM	o1F]��O\�y\JDaИ#�x���f�)�'a
�M~�L~:?�׾���'?�&?Kko	no	VZ��VD�YB?BL��e��	!�o��t��H|�Mv���Ӿ/na'~n!2Hke�nM�Vp��f]�y?jDYLH�!S��a�g�8�&��OM~�#i|�o�Ӿ���%3�'>VZO	o
�V\�VL�AJNY@`!S��6�=S2k�n��h��Dh��ea��Eql�T�VQoZ_��f��fmc�,aCc�MW@Wc�ҽf�7g,�WE�ʽ�½2�o��j���h��ws��Es��T}�SPC[��d�C�byC��mA�' ,a�©6ƬrO�j_.�b�lh��Es�Ew��P?�g��	�f��&lC�iO�$3L �f��7�A.3O��A��h�lE`�Er�}�~�}Pz�0�f��viC�,`A�,(G1�5=�µO(7{S-�h��hlTs��Wc��@o�_@�O��f4�faSk�iC� �BBY�B=[SO�O��`��&h��%sx-%`��pp�P;�V�+�"4�fqC�a[�<	Q�&¿��2K� C��`�d�(�heq}KWs�py�_@�X�+f��&iC��h�,!$���6�?M�J*�h��x��es}�rw�ER�KR~S{�d�/�fqg�iA� 5U�½&�_�[��h�n�j��%3l�er��P}�oSuYOu
_b\�li�hC�,@6F�6��O�O��i�h dEa��Ar�OP��]Xm�^�	�f��fHC�,)a+�,A������33G�O��h��h��Es�Mas�@�Vw}_�+~l�
�faF�,iCg<AI�b��¼^�O�& ��h��Es݇c��P?�_@oKW0V�d��mi��iCk�tA
ݶ�%0��J��c�lFh�p�/As��PJUP�}��g�	�b(c)�mC��3%a���6.B10SO�0R[.�h��x��Es}�ec�-P{XmsW�C�f��gmC��hC�D7 ���:
�RCO�N��(��x�as��Es}p�]P_�N��j��fi�ic� :�r;g�d�$N*Y%Ff�M"�M��: s�:*��*������*��|m�Pty� "��"�1�{ggd*�`
�$
�,nj�M�b�m��:��r ��ڪ�,���V��*4�ph�uh�"��"�(��"�E&th�th�".�"�3�)�t;g�l
�:N
I$Nf�-Ob�Ms�(Ps�:k�X�[*����4�tdt`� "�2�2�;ge/���lK
�$Nb�	�b���d8 ��:�n��*��B�j��k4�ph4tl�"�� �1 *o�l?�d�$L�dOb�Lg�����2��Z�렚�b�*��th�tl["��b��+��l;��d�&N
�$jbPMb������:��آ��Ҩ�����qh�phSP".�"��;�l;�d�$ �$nb�%} �?]q�:p��:�k�Z���گ�4�j��dh�0`�!b�W"��8|� ;o�d
I&NB4Nf�'�b���*0��:P�{�z��,ڪ�����el�p)�"��"��Ee?�d
�$N
I�Ff�]C�-��D;��sd*�ڠ��"����u`�v`�#�� ��dkgpI4J�,Nb�6�hT���:Q�D;"k��Z�$ڨ� ���\�th�  (� ",�b��+�g9�d�&N
�4Nj�-�b���:��*@(�l�*��j�*�bvh0d(�5ݮ"��;�d)�t�$j�$L@��c�	�s�FUqT9"�J�˄ڪ����"th�0th+";"� uG�d+�:� F� ^r��bTM��:��:)�X���Һ�����th�t}�0&�1�.�{�l+�t:�dNr�$^b�LDN�M���{0s�( 
�˫{�Ī�����5(vy� ��".�:�f?�FD�&NB�$Nb�M�j�E�p2��20*�r��ڢ(���"t(�dh�#��"��Mb��]��`�O���/b��