.1�
/1--},-}.,!7I)1M/�e/z	e<s9??�41v�<8��pI��`I��,��L#.3
.� -}*�}
!7KD!3K.jK�/�K�2sV8sv�5p~�4d�� 	��`M��
%��.1�	.��-}.�}%7I%3O/zm/:e<383-�51~�40��`i��!i��
����*#� .1E@�t*(!uBLa3K! K�e/z�!w0sFv�4xw�<0��tI�� ����#.3�,���}*-}*%5K!3-��-�m<s8sd�44w�,0��0I��pI�F#��'/�%,1�B-uF-}ZH+2J)O+Zm/�e/s8sv�<0t�48�� i��1M��%��#/#%-�-�=�}*-)3O)3K-�-�e8'8su�40V�4p��pK��`i�B#��.�� .�-}(�m*,)7!?K/�e/>	�8c8su�4,w�48��`I��`I������.�..%��},�}+,!K3/Ze*�c839{g�4%v�4%��0m��ti�#��.��.��-}
-m/,!!O$!3K/��/�	�91<q/�54o�< ��bm��qi��R!��X",��.���u"�,
l 3KD)3O�Ce+�E0sF8st�|<v�>q��li��hi�FZ#�FZ!.��R)#�B)}*,�x,%6[ #K?�e's/�8w4,Vr�4tr�40��pi��`I�LO���#+7�F.�%�t
$)}J-3J!2O@/�e_r	�W8qV?8aFg�18r�t ��rH��pi��^#�F�.�B.3�!-d*h-x*!0J!#I/~g-��8u8uVv�<0f�48��pi��`i�Nb�F�(�� .:��mkL-}o!;Z)#[�Cu/�A�<c8s[r�/0v�4t��rI��0	��!��!.3�&3�B�|*,%}Ho%sKDa3AD.xOe?�e:sUxsT��40v�|p��bA��pM�D^#���$��T)ak|cil��Ar��Or�3�N1�%؍i�܁<ae-aE"aV�r�v�@^�P@��_5$$^D`�o/�C�iL��Kr��Kv�5�N"�)���i�܉nQElcD"C_�g�v�P��DN��.$��h��k�#bKlC��b��Cb�;��q�(��-&ށlcv,ce#Kt�&K^�@-�X@V���t$$^ ��a,B�k���r��#j�3�V3�m$͉)��	)ce_(Ce]f{R� �U�DL��E���"�� 4�h�#ci�*��Cr��AxN3�^;�a��)m�$cEM(se2KU�b�w�@!�p@��V 4^$��il�k�#��r��p�'��s�m�܈+�č,`E]dsE&Kv�bkv�L�hH�/�4 0^1��)?#�i���~��bL;��;�)݉)��	,cE,cE&k�"k>�I�m@��^$�O4 �c-�#oml#��z��b+��3�)��	)���laF$re"mu�2KW�@�Q@�P�.t_(��)lcjh��r��p^g�V1�i/�Ii܉8/E-cDMf�^�*�v�@��@��.u`4� �ky�#�i�2��Cb��Cb�#��2�)&܁s�	Se,ba]"�~�"kV�B��@�H^ 4^T �Kh# ���w��b^?�R7�)�	)�SE]KGO"z4�&Ku�@��P�P�"�V4b2ci(�h���q��p#�Z3�?!2܉I���lca,bErK^�b*6�@�P �@^p4�U`fcimcih��r��rJ#�2�_+�	l�܍mcI:BE �V�2kV�@
�p@�`�T �^t ��kf#�i���r��s^2��2�)n܉)��mkE_,cE"�t�"[V�@^��@��Z4���4a�cyl�il#��p��CbR?�\3�)���n�ܙlgM-gIc�V�"�V�A�P@�PD-��5 �cl�i`��r��r��n��|)3`+1`[4��I51��T�|�tO� E�@P]W[�#K4���4N9�v�| Eo:OwV�"��#�&._.�_�Qd�e1n�������)03`-)3`A0 �Cp2��t�2�uV� �rEwd�#��1�&�_�_�qt��1`������� Y3biY3`0��4���t�>�dL�@-vRPDwP�"��&�&�Kf�O�uf��1d���N��\)3(){`Kt��
4���T�:�T�xE�ZCgt�#��!�"�_.�_gt�cqd���\���HU1c)3`Ku0�m4 ��4θ�t�t!sR Ewb�3��+�&�N �_ful��q`���~���+3`)3dKt��C$���T��T_8oczef1�"��!� '�_&�Kg1h�#3d���N���9	3 	YsdKt��K>���vO<�uN�EwR GgR�#��#�n�"�AW�; �'1d�������)3d!93`Kv��K4���t8�p8UWRMwR�g�&�3�&�H6�Ocs`�#1d���^��^	3p)sck-0�K$0��t���@8 E�V DgR1#��'�*�&�f1d��1d�N���N���%93 9h7b4 �0 ��F��t@� EwREgr�#��#�&�&�^e0 �g1d������~l3`)9#aJt�K4���TN8�tN�A�b@/p�"��#�	&�AI"�N�3d��se���~���)# )13`i0 �Z4���T��TθE7RE�X�#��#�$� W&�Ogqe��d�����* 9#`)93  $0�C5���eN��T^� �r U�r� ��#�'�Vf�O�q`�oud������n)93`+#hYt��Kv0��t�4�TN�$fAsP�//�#�&�_$�^a1d��1 �������)3*)93 C4��i=���4J8�T�8 DbrHE�s�#� �!� �].� O�9 �g1`����=}��u,�1)�d1�ea��`% !�% !⮝ i��!�:Ց�8���i�������8�������}���1)�d5)�$g�U)�}��-w��-5)�d})(�g��av��ob(�E #��� y�� ���롸�Щ��������
����u�=|��w5+��=)��w�WgW��kE:+�  �� q�� �����������������0�>���}��}��1),�1(,�w��kv�Uc%=r )r�� �� !+���8���p������������}��45)v�5!��w��k5�/k!	� !�� �� �:Ǔ��������ñ�8��: ���m��}�ε%(��4)�df��kg�U{%$)�%)������ .����8���i�������0���>i��=m���4)�d1)l�'�E+�Di! !� (`�� � 񺦲�8�������x���p��:0�Ֆ�����=5)�au)�fw�ui6�Eb )r (2��y��@�𷓩8���h���������<������<|��1(�d1)9�W�Ugw�+@Hr i�� ��� �4ד�9�����������<���0��^���=���%(l�5)l�w�Ukw��kA)r%*)