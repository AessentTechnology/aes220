----------------------------------------------------------------------------------------------------
-- File name: AsymmetricS16S16DualPortRAM_V1.0.0.vhd
----------------------------------------------------------------------------------------------------
-- Author: Sebastien Saury, Aessent Technology Ltd
----------------------------------------------------------------------------------------------------
-- DESCRIPTION
--
-- Instantiates a BRAM with a 16 bit port on both sides
-- No parity signal used. 
--
----------------------------------------------------------------------------------------------------
--CHANGES
--
-- V1.0.0: original version
-- 
----------------------------------------------------------------------------------------------------
--NOTES
--
-- Original template from RAMB16_S18_S9 comes from Xilinx own documentation
--
----------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2012-2013 Sebastien Saury, Aessent Technology Ltd
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the Lesser GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
----------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;             -- Required for BRAM instantiation

entity S16S16_dual_port_RAM_ent is

  port (
    CLKA_in  : in  std_logic;
    CLKB_in  : in  std_logic;
    ENA_in   : in  std_logic;
    ENB_in   : in  std_logic;
    WEA_in   : in  unsigned(1 downto 0);
    WEB_in   : in  std_logic;
    ADDRA_in : in  unsigned(9 downto 0);
    ADDRB_in : in  unsigned(9 downto 0);
    DIA_in   : in  unsigned(15 downto 0);
    DIB_in   : in  unsigned(15 downto 0);
    DOA_out  : out unsigned(15 downto 0);
    DOB_out  : out unsigned(15 downto 0));

end S16S16_dual_port_RAM_ent;

architecture instantiation_arch of S16S16_dual_port_RAM_ent is

  signal doa_s : std_logic_vector(15 downto 0);
  signal dob_s : std_logic_vector(15 downto 0);

begin

   -- RAMB16_S18_S9: 1k/2k x 16/8 + 2/1 Parity bit Dual-Port RAM
   --               Spartan-3A
   -- Xilinx HDL Language Template, version 14.2

   RAMB16_S16S16_inst : RAMB16BWE_S18_S18
   generic map (
      INIT_A => x"00000", --  Value of output RAM registers on Port A at startup
      INIT_B => x"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => x"00000", --  Port A output value upon SSR assertion
      SRVAL_B => x"00000", --  Port B output value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL"
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Port A Address 0 to 255, Port B Address 0 to 255
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 256 to 511, Port B Address 256 to 511
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 512 to 767, Port B Address 1024 to 1535
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 768 to 1023, Port B Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      CLKA => CLKA_in,    -- Port A Clock
      CLKB => CLKB_in,    -- Port B Clock
      ENA => ENA_in,      -- Port A RAM Enable Input
      ENB => ENB_in,      -- PortB RAM Enable Input
      SSRA => '0',        -- Port A Synchronous Set/Reset Input
      SSRB => '0',        -- Port B Synchronous Set/Reset Input
      WEA => std_logic_vector(WEB_in),     -- Port A 2-bit Write Enable Input
      WEB => std_logic_vector(WEB_in),     -- Port B 2-bit Write Enable Input
      ADDRA => std_logic_vector(ADDR_in),  -- Port A 11-bit Address Input
      ADDRB => std_logic_vector(ADDR_in),  -- Port B 11-bit Address Input
      DIA => std_logic_vector(DIA_in),     -- Port A 16-bit Data Input
      DIB => std_logic_vector(DIB_in),     -- Port B 16-bit Data Input
      DIPA => "00",        -- Port A 2-bit parity
      DIPB => "00",        -- Port B 2-bit parity
      DOA => doa_s,     -- Port A 16-bit Data Output
      DOB => dob_s);    -- Port B 16-bit Data Output

   DOA_out <= unsigned(doa_s);
   DOB_out <= unsigned(dob_s);
  
end instantiation_arch;
